-- Code your testbench here
library IEEE;
use IEEE.std_logic_1164.all;

entity TOP_TMR is
end TOP_TMR;

architecture TMR_ARCHITECTURE of TOP_TMR is

component TMR is
port (	
  i_CANAL1 	:  in std_logic_vector(15 downto 0); -- Entrada 1 de dados
  i_CANAL2 	:  in std_logic_vector(15 downto 0); -- Entrada 2 de dados
  i_CANAL3 	:  in std_logic_vector(15 downto 0); -- Entrada 3 de dados
  o_RETURN  :  out std_logic_vector(15 downto 0)); -- Saida de dados
end component;

signal w_END: std_logic_vector (15 downto 0);-- Definir signal w_END
signal w_S: std_logic_vector (15 downto 0); -- Definir signal w_S
signal w_1: std_logic_vector (15 downto 0); -- Definir signal w_1
signal w_2: std_logic_vector (15 downto 0); -- Definir signal w_2
signal w_3: std_logic_vector (15 downto 0); -- Definir signal w_3

begin
u_TMR: TMR port map( -- Definir as portas do TMR
  i_CANAL1  =>  w_1,
  i_CANAL2  =>  w_2,
  i_CANAL3  =>  w_3,
  o_RETURN  =>  w_S);

process
begin
-- Primeiro teste para checar se a função do VOTER esta certo para i_1 == i_2
w_1  <=  "1010101010101010";
w_2  <=  "1010101010101010";
w_3	 <=  "1010101010101011";
wait for 3ns;
assert (w_S  =  "0000000000000000") report "Falha no teste 1" severity error;

-- Segundo teste para checar se a função do VOTER esta certo para i_1 == i_3
w_1  <=  "1100110011001100";
w_2  <=  "0011110000111100";
w_3	 <=  "1100110011001100";
wait for 3ns;
assert (w_S  =  "0000000000000000") report "Falha no teste 2" severity error;

-- Terceiro teste para chegar se a função do VOTER esta certo para i_2 == i_3
w_1 <= "1111111111111111";
w_2 <= "0000000011111111";
w_3	<= "0000000011111111";
wait for 3ns;
assert (w_S  =  "0000000000000000") report "Falha no teste 3" severity error;

-- Quarto teste para chegar se a função do VOTER esta certo para i_1 == i_2 == i_3
w_1 <= "0000000011111111";
w_2 <= "0000000011111111";
w_3	<= "0000000011111111";
wait for 3ns;
assert (w_S  =  "0000000000000000") report "Falha no teste 4" severity error;

-- Limpar os dados w_1, w_2 e w_3
      w_1  <=  "0000000000000000";
      w_2  <=  "0000000000000000";
      w_3  <=  "0000000000000000";
      wait for 1ns;
      assert false report "Teste Concluido." severity note; --Avisa se o teste teve exito
      end process;
      end architecture;